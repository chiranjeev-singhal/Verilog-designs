module decimal ();

reg [2:0] deci;

initial
begin
deci = 3'd4;
$display (deci);
end
endmodule 
